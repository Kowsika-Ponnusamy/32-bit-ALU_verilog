module prefix32pipe(s,cout,a,b,c,clk,reset);
input [31:0] a,b;
input c,clk,reset;
output[31:0] s;
output cout;
wire [31:0] p,g,k;
wire [31:0] x;
wire [63:0] df0;
wire [61:0] df1;
wire [57:0] df2;
wire [49:0] df3;
wire [33:0] df4,df5;
wire cout1,cout2;
assign p=a^b;
assign g=a&b;
assign k=g|p;
wire g12,g34,g56,g78,g910,g1112,g1314,g1516,g1718,g1920,g2122,g2324,g2526,g2728,g2930,g35,g36,g79,g710,g711,g712,g713,g714,g1113,g1114,g1921,g1922,g2325,g2326,g2729,g2730;
wire k12,k34,k56,k78,k910,k1112,k1314,k1516,k1718,k1920,k2122,k2324,k2526,k2728,k2930,k35,k36,k79,k710,k711,k712,k713,k714,k1113,k1114,k1921,k1922,k2325,k2326,k2729,k2730;
wire g1517,g1518,g1519,g1520,g1521,g1522,g1523,g1524,g1525,g1526,g1527,g1528,g1529,g1530,g2327,g2328,g2329,g2330;
wire k1517,k1518,k1519,k1520,k1521,k1522,k1523,k1534,k1525,k1526,k1527,k1528,k1529,k1530,k2327,k2328,k2329,k2330;
assign x[0]=c;
//stage 1
dot d1(x[1],g[0],k[0],x[0]);
circle c1(g[2],k[2],g[1],k[1],g12,k12);
circle c2(g[4],k[4],g[3],k[3],g34,k34);
circle c3(g[6],k[6],g[5],k[5],g56,k56);
circle c4(g[8],k[8],g[7],k[7],g78,k78);
circle c5(g[10],k[10],g[9],k[9],g910,k910);
circle c6(g[12],k[12],g[11],k[11],g1112,k1112);
circle c7(g[14],k[14],g[13],k[13],g1314,k1314);
circle c8(g[16],k[16],g[15],k[15],g1516,k1516);
circle c9(g[18],k[18],g[17],k[17],g1718,k1718);
circle c10(g[20],k[20],g[19],k[19],g1920,k1920);
circle c11(g[22],k[22],g[21],k[21],g2122,k2122);
circle c12(g[24],k[24],g[23],k[23],g2324,k2324);
circle c13(g[26],k[26],g[25],k[25],g2526,k2526);
circle c14(g[28],k[28],g[27],k[27],g2728,k2728);
circle c15(g[30],k[30],g[29],k[29],g2930,k2930);
d_ff dff000(x[0],clk,reset,df0[0]);
d_ff dff001(x[1],clk,reset,df0[1]);
d_ff dff002(g[1],clk,reset,df0[2]);
d_ff dff003(k[1],clk,reset,df0[3]);
d_ff dff004(g12,clk,reset,df0[4]);
d_ff dff005(k12,clk,reset,df0[5]);
d_ff dff006(g[3],clk,reset,df0[6]);
d_ff dff007(k[3],clk,reset,df0[7]);
d_ff dff008(g34,clk,reset,df0[8]);
d_ff dff009(k34,clk,reset,df0[9]);
d_ff dff010(g[5],clk,reset,df0[10]);
d_ff dff011(k[5],clk,reset,df0[11]);
d_ff dff012(g56,clk,reset,df0[12]);
d_ff dff013(k56,clk,reset,df0[13]);
d_ff dff014(g[7],clk,reset,df0[14]);
d_ff dff015(k[7],clk,reset,df0[15]);
d_ff dff016(g78,clk,reset,df0[16]);
d_ff dff017(k78,clk,reset,df0[17]);
d_ff dff018(g[9],clk,reset,df0[18]);
d_ff dff019(k[9],clk,reset,df0[19]);
d_ff dff020(g910,clk,reset,df0[20]);
d_ff dff021(k910,clk,reset,df0[21]);
d_ff dff022(g[11],clk,reset,df0[22]);
d_ff dff023(k[11],clk,reset,df0[23]);
d_ff dff024(g1112,clk,reset,df0[24]);
d_ff dff025(k1112,clk,reset,df0[25]);
d_ff dff026(g[13],clk,reset,df0[26]);
d_ff dff027(k[13],clk,reset,df0[27]);
d_ff dff028(g1314,clk,reset,df0[28]);
d_ff dff029(k1314,clk,reset,df0[29]);
d_ff dff030(g[15],clk,reset,df0[30]);
d_ff dff031(k[15],clk,reset,df0[31]);
d_ff dff032(g1516,clk,reset,df0[32]);
d_ff dff033(k1516,clk,reset,df0[33]);
d_ff dff034(g[17],clk,reset,df0[34]);
d_ff dff035(k[17],clk,reset,df0[35]);
d_ff dff036(g1718,clk,reset,df0[36]);
d_ff dff037(k1718,clk,reset,df0[37]);
d_ff dff038(g[19],clk,reset,df0[38]);
d_ff dff039(k[19],clk,reset,df0[39]);
d_ff dff040(g1920,clk,reset,df0[40]);
d_ff dff041(k1920,clk,reset,df0[41]);
d_ff dff042(g[21],clk,reset,df0[42]);
d_ff dff043(k[21],clk,reset,df0[43]);
d_ff dff044(g2122,clk,reset,df0[44]);
d_ff dff045(k2122,clk,reset,df0[45]);
d_ff dff046(g[23],clk,reset,df0[46]);
d_ff dff047(k[23],clk,reset,df0[47]);
d_ff dff048(g2324,clk,reset,df0[48]);
d_ff dff049(k2324,clk,reset,df0[49]);
d_ff dff050(g[25],clk,reset,df0[50]);
d_ff dff051(k[25],clk,reset,df0[51]);
d_ff dff052(g2526,clk,reset,df0[52]);
d_ff dff053(k2526,clk,reset,df0[53]);
d_ff dff054(g[27],clk,reset,df0[54]);
d_ff dff055(k[27],clk,reset,df0[55]);
d_ff dff056(g2728,clk,reset,df0[56]);
d_ff dff057(k2728,clk,reset,df0[57]);
d_ff dff058(g[29],clk,reset,df0[58]);
d_ff dff059(k[29],clk,reset,df0[59]);
d_ff dff060(g2930,clk,reset,df0[60]);
d_ff dff061(k2930,clk,reset,df0[61]);
d_ff dff062(g[31],clk,reset,df0[62]);
d_ff dff063(k[31],clk,reset,df0[63]);
//stage 2
dot d2(x[2],df0[2],df0[3],df0[1]);
dot d3(x[3],df0[4],df0[5],df0[1]);
circle c16(df0[10],df0[11],df0[8],df0[9],g35,k35);
circle c17(df0[12],df0[13],df0[8],df0[9],g36,k36);
circle c18(df0[18],df0[19],df0[16],df0[17],g79,k79);
circle c19(df0[20],df0[21],df0[16],df0[17],g710,k710);
circle c20(df0[26],df0[27],df0[24],df0[25],g1113,k1113);
circle c21(df0[28],df0[29],df0[24],df0[25],g1114,k1114);
circle c22(df0[34],df0[35],df0[32],df0[33],g1517,k1517);
circle c23(df0[36],df0[37],df0[32],df0[33],g1518,k1518);
circle c24(df0[42],df0[43],df0[40],df0[41],g1921,k1921);
circle c25(df0[44],df0[45],df0[40],df0[41],g1922,k1922);
circle c26(df0[50],df0[51],df0[48],df0[49],g2325,k2325);
circle c27(df0[52],df0[53],df0[48],df0[49],g2326,k2326);
circle c28(df0[58],df0[59],df0[56],df0[57],g2729,k2729);
circle c29(df0[60],df0[61],df0[56],df0[57],g2730,k2730);
d_ff dff100(df0[0],clk,reset,df1[0]);
d_ff dff101(df0[1],clk,reset,df1[1]);
d_ff dff102(x[2],clk,reset,df1[2]);
d_ff dff103(x[3],clk,reset,df1[3]);
d_ff dff104(df0[6],clk,reset,df1[4]);
d_ff dff105(df0[7],clk,reset,df1[5]);
d_ff dff106(df0[8],clk,reset,df1[6]);
d_ff dff107(df0[9],clk,reset,df1[7]);
d_ff dff108(g35,clk,reset,df1[8]);
d_ff dff109(k35,clk,reset,df1[9]);
d_ff dff110(g36,clk,reset,df1[10]);
d_ff dff111(k36,clk,reset,df1[11]);
d_ff dff112(df0[14],clk,reset,df1[12]);
d_ff dff113(df0[15],clk,reset,df1[13]);
d_ff dff114(df0[16],clk,reset,df1[14]);
d_ff dff115(df0[17],clk,reset,df1[15]);
d_ff dff116(g79,clk,reset,df1[16]);
d_ff dff117(k79,clk,reset,df1[17]);
d_ff dff118(g710,clk,reset,df1[18]);
d_ff dff119(k710,clk,reset,df1[19]);
d_ff dff120(df0[22],clk,reset,df1[20]);
d_ff dff121(df0[23],clk,reset,df1[21]);
d_ff dff122(df0[24],clk,reset,df1[22]);
d_ff dff123(df0[25],clk,reset,df1[23]);
d_ff dff124(g1113,clk,reset,df1[24]);
d_ff dff125(k1113,clk,reset,df1[25]);
d_ff dff126(g1114,clk,reset,df1[26]);
d_ff dff127(k1114,clk,reset,df1[27]);
d_ff dff128(df0[30],clk,reset,df1[28]);
d_ff dff129(df0[31],clk,reset,df1[29]);
d_ff dff130(df0[32],clk,reset,df1[30]);
d_ff dff131(df0[33],clk,reset,df1[31]);
d_ff dff132(g1517,clk,reset,df1[32]);
d_ff dff133(k1517,clk,reset,df1[33]);
d_ff dff134(g1518,clk,reset,df1[34]);
d_ff dff135(k1518,clk,reset,df1[35]);
d_ff dff136(df0[38],clk,reset,df1[36]);
d_ff dff137(df0[39],clk,reset,df1[37]);
d_ff dff138(df0[40],clk,reset,df1[38]);
d_ff dff139(df0[41],clk,reset,df1[39]);
d_ff dff140(g1921,clk,reset,df1[40]);
d_ff dff141(k1921,clk,reset,df1[41]);
d_ff dff142(g1922,clk,reset,df1[42]);
d_ff dff143(k1922,clk,reset,df1[43]);
d_ff dff144(df0[46],clk,reset,df1[44]);
d_ff dff145(df0[47],clk,reset,df1[45]);
d_ff dff146(df0[48],clk,reset,df1[46]);
d_ff dff147(df0[49],clk,reset,df1[47]);
d_ff dff148(g2325,clk,reset,df1[48]);
d_ff dff149(k2325,clk,reset,df1[49]);
d_ff dff150(g2326,clk,reset,df1[50]);
d_ff dff151(k2326,clk,reset,df1[51]);
d_ff dff152(df0[54],clk,reset,df1[52]);
d_ff dff153(df0[55],clk,reset,df1[53]);
d_ff dff154(df0[56],clk,reset,df1[54]);
d_ff dff155(df0[57],clk,reset,df1[55]);
d_ff dff156(g2729,clk,reset,df1[56]);
d_ff dff157(k2729,clk,reset,df1[57]);
d_ff dff158(g2730,clk,reset,df1[58]);
d_ff dff159(k2730,clk,reset,df1[59]);
d_ff dff160(df0[60],clk,reset,df1[60]);
d_ff dff161(df0[61],clk,reset,df1[61]);
//stage 3

dot d4(x[4],df1[4],df1[5],df1[3]);
dot d5(x[5],df1[6],df1[7],df1[3]);
dot d6(x[6],df1[8],df1[9],df1[3]);
dot d7(x[7],df1[10],df1[11],df1[3]);
circle c30(df1[20],df1[21],df1[18],df1[19],g711,k711);
circle c31(df1[22],df1[23],df1[18],df1[19],g712,k712);
circle c32(df1[24],df1[25],df1[18],df1[19],g713,k713);
circle c33(df1[26],df1[27],df1[18],df1[19],g714,k714);
circle c34(df1[36],df1[37],df1[34],df1[35],g1519,k1519);
circle c35(df1[38],df1[39],df1[34],df1[35],g1520,k1520);
circle c36(df1[40],df1[41],df1[34],df1[35],g1521,k1521);
circle c37(df1[42],df1[43],df1[34],df1[35],g1522,k1522);
circle c38(df1[52],df1[53],df1[50],df1[51],g2327,k2327);
circle c39(df1[54],df0[55],df1[50],df1[51],g2328,k2328);
circle c40(df1[56],df1[57],df1[50],df1[51],g2329,k2329);
circle c41(df1[58],df1[59],df1[50],df1[51],g2330,k2330);
d_ff dff200(df1[0],clk,reset,df2[0]);
d_ff dff201(df1[1],clk,reset,df2[1]);
d_ff dff202(df1[2],clk,reset,df2[2]);
d_ff dff203(df1[3],clk,reset,df2[3]);
d_ff dff204(x[4],clk,reset,df2[4]);
d_ff dff205(x[5],clk,reset,df2[5]);
d_ff dff206(x[6],clk,reset,df2[6]);
d_ff dff207(x[7],clk,reset,df2[7]);
d_ff dff208(df1[12],clk,reset,df2[8]);
d_ff dff209(df1[13],clk,reset,df2[9]);
d_ff dff210(df1[14],clk,reset,df2[10]);
d_ff dff211(df1[15],clk,reset,df2[11]);
d_ff dff212(df1[16],clk,reset,df2[12]);
d_ff dff213(df1[17],clk,reset,df2[13]);
d_ff dff214(df1[18],clk,reset,df2[14]);
d_ff dff215(df1[19],clk,reset,df2[15]);
d_ff dff216(g711,clk,reset,df2[16]);
d_ff dff217(k711,clk,reset,df2[17]);
d_ff dff218(g712,clk,reset,df2[18]);
d_ff dff219(k712,clk,reset,df2[19]);
d_ff dff220(g713,clk,reset,df2[20]);
d_ff dff221(k713,clk,reset,df2[21]);
d_ff dff222(g714,clk,reset,df2[22]);
d_ff dff223(k714,clk,reset,df2[23]);
d_ff dff224(df1[28],clk,reset,df2[24]);
d_ff dff225(df1[29],clk,reset,df2[25]);
d_ff dff226(df1[30],clk,reset,df2[26]);
d_ff dff227(df1[31],clk,reset,df2[27]);
d_ff dff228(df1[32],clk,reset,df2[28]);
d_ff dff229(df1[33],clk,reset,df2[29]);
d_ff dff230(df1[34],clk,reset,df2[30]);
d_ff dff231(df1[35],clk,reset,df2[31]);
d_ff dff232(g1519,clk,reset,df2[32]);
d_ff dff233(k1519,clk,reset,df2[33]);
d_ff dff234(g1520,clk,reset,df2[34]);
d_ff dff235(k1520,clk,reset,df2[35]);
d_ff dff236(g1521,clk,reset,df2[36]);
d_ff dff237(k1521,clk,reset,df2[37]);
d_ff dff238(g1522,clk,reset,df2[38]);
d_ff dff239(k1522,clk,reset,df2[39]);
d_ff dff240(df1[44],clk,reset,df2[40]);
d_ff dff241(df1[45],clk,reset,df2[41]);
d_ff dff242(df1[46],clk,reset,df2[42]);
d_ff dff243(df1[47],clk,reset,df2[43]);
d_ff dff244(df1[48],clk,reset,df2[44]);
d_ff dff245(df1[49],clk,reset,df2[45]);
d_ff dff246(df1[50],clk,reset,df2[46]);
d_ff dff247(df1[51],clk,reset,df2[47]);
d_ff dff248(g2327,clk,reset,df2[48]);
d_ff dff249(k2327,clk,reset,df2[49]);
d_ff dff250(g2328,clk,reset,df2[50]);
d_ff dff251(k2328,clk,reset,df2[51]);
d_ff dff252(g2329,clk,reset,df2[52]);
d_ff dff253(k2329,clk,reset,df2[53]);
d_ff dff254(g2330,clk,reset,df2[54]);
d_ff dff255(k2330,clk,reset,df2[55]);
d_ff dff256(df1[60],clk,reset,df2[56]);
d_ff dff257(df1[61],clk,reset,df2[57]);
//stage 4
dot d8(x[8],df2[8],df2[9],df2[7]);
dot d9(x[9],df2[10],df2[11],df2[7]);
dot d10(x[10],df2[12],df2[13],df2[7]);
dot d11(x[11],df2[14],df1[15],df2[7]);
dot d12(x[12],df2[16],df2[17],df2[7]);
dot d13(x[13],df2[18],df2[19],df2[7]);
dot d14(x[14],df2[20],df2[21],df2[7]);
dot d15(x[15],df2[22],df2[23],df2[7]);
circle c42(df2[40],df2[41],df2[38],df2[39],g1523,k1523);
circle c43(df2[42],df2[43],df2[38],df2[39],g1524,k1524);
circle c44(df2[44],df2[45],df2[38],df2[39],g1525,k1525);
circle c45(df2[46],df2[47],df2[38],df2[39],g1526,k1526);
circle c46(df2[48],df2[49],df2[38],df2[39],g1527,k1527);
circle c47(df2[50],df2[51],df2[38],df2[39],g1528,k1528);
circle c48(df2[52],df2[53],df2[38],df2[39],g1529,k1529);
circle c49(df2[54],df2[55],df2[38],df2[39],g1530,k1530);
d_ff dff300(df2[0],clk,reset,df3[0]);
d_ff dff301(df2[1],clk,reset,df3[1]);
d_ff dff302(df2[2],clk,reset,df3[2]);
d_ff dff303(df2[3],clk,reset,df3[3]);
d_ff dff304(df2[4],clk,reset,df3[4]);
d_ff dff305(df2[5],clk,reset,df3[5]);
d_ff dff306(df2[6],clk,reset,df3[6]);
d_ff dff307(df2[7],clk,reset,df3[7]);
d_ff dff308(x[8],clk,reset,df3[8]);
d_ff dff309(x[9],clk,reset,df3[9]);
d_ff dff310(x[10],clk,reset,df3[10]);
d_ff dff311(x[11],clk,reset,df3[11]);
d_ff dff312(x[12],clk,reset,df3[12]);
d_ff dff313(x[13],clk,reset,df3[13]);
d_ff dff314(x[14],clk,reset,df3[14]);
d_ff dff315(x[15],clk,reset,df3[15]);
d_ff dff316(df2[24],clk,reset,df3[16]);
d_ff dff317(df2[25],clk,reset,df3[17]);
d_ff dff318(df2[26],clk,reset,df3[18]);
d_ff dff319(df2[27],clk,reset,df3[19]);
d_ff dff320(df2[28],clk,reset,df3[20]);
d_ff dff321(df2[29],clk,reset,df3[21]);
d_ff dff322(df2[30],clk,reset,df3[22]);
d_ff dff323(df2[31],clk,reset,df3[23]);
d_ff dff324(df2[32],clk,reset,df3[24]);
d_ff dff325(df2[33],clk,reset,df3[25]);
d_ff dff326(df2[34],clk,reset,df3[26]);
d_ff dff327(df2[35],clk,reset,df3[27]);
d_ff dff328(df2[36],clk,reset,df3[28]);
d_ff dff329(df2[37],clk,reset,df3[29]);
d_ff dff330(df2[38],clk,reset,df3[30]);
d_ff dff331(df2[39],clk,reset,df3[31]);
d_ff dff332(g1523,clk,reset,df3[32]);
d_ff dff333(k1523,clk,reset,df3[33]);
d_ff dff334(g1524,clk,reset,df3[34]);
d_ff dff335(k1524,clk,reset,df3[35]);
d_ff dff336(g1525,clk,reset,df3[36]);
d_ff dff337(k1525,clk,reset,df3[37]);
d_ff dff338(g1526,clk,reset,df3[38]);
d_ff dff339(k1526,clk,reset,df3[39]);
d_ff dff340(g1527,clk,reset,df3[40]);
d_ff dff341(k1527,clk,reset,df3[41]);
d_ff dff342(g1528,clk,reset,df3[42]);
d_ff dff343(k1528,clk,reset,df3[43]);
d_ff dff344(g1529,clk,reset,df3[44]);
d_ff dff345(k1529,clk,reset,df3[45]);
d_ff dff346(g1530,clk,reset,df3[46]);
d_ff dff347(k1530,clk,reset,df3[47]);
d_ff dff348(df2[56],clk,reset,df3[48]);
d_ff dff349(df2[57],clk,reset,df3[49]);
//stage 5
dot d16(x[16],df3[16],df3[17],df3[15]);
dot d17(x[17],df3[18],df3[19],df3[15]);
dot d18(x[18],df3[20],df3[21],df3[15]);
dot d19(x[19],df3[22],df3[23],df3[15]);
dot d20(x[20],df3[24],df3[25],df3[15]);
dot d21(x[21],df3[26],df3[27],df3[15]);
dot d22(x[22],df3[28],df3[29],df3[15]);
dot d23(x[23],df3[30],df3[31],df3[15]);
dot d24(x[24],df3[32],df3[33],df3[15]);
dot d25(x[25],df3[34],df3[35],df3[15]);
dot d26(x[26],df3[36],df3[37],df3[15]);
dot d27(x[27],df3[38],df3[39],df3[15]);
dot d28(x[28],df3[40],df3[41],df3[15]);
dot d29(x[29],df3[42],df3[43],df3[15]);
dot d30(x[30],df3[44],df3[45],df3[15]);
dot d31(x[31],df3[46],df3[47],df3[15]);
d_ff dff400(df3[0],clk,reset,df4[0]);
d_ff dff401(df3[1],clk,reset,df4[1]);
d_ff dff402(df3[2],clk,reset,df4[2]);
d_ff dff403(df3[3],clk,reset,df4[3]);
d_ff dff404(df3[4],clk,reset,df4[4]);
d_ff dff405(df3[5],clk,reset,df4[5]);
d_ff dff406(df3[6],clk,reset,df4[6]);
d_ff dff407(df3[7],clk,reset,df4[7]);
d_ff dff408(df3[8],clk,reset,df4[8]);
d_ff dff409(df3[9],clk,reset,df4[9]);
d_ff dff410(df3[10],clk,reset,df4[10]);
d_ff dff411(df3[11],clk,reset,df4[11]);
d_ff dff412(df3[12],clk,reset,df4[12]);
d_ff dff413(df3[13],clk,reset,df4[13]);
d_ff dff414(df3[14],clk,reset,df4[14]);
d_ff dff415(df3[15],clk,reset,df4[15]);
d_ff dff416(x[16],clk,reset,df4[16]);
d_ff dff417(x[17],clk,reset,df4[17]);
d_ff dff418(x[18],clk,reset,df4[18]);
d_ff dff419(x[19],clk,reset,df4[19]);
d_ff dff420(x[20],clk,reset,df4[20]);
d_ff dff421(x[21],clk,reset,df4[21]);
d_ff dff422(x[22],clk,reset,df4[22]);
d_ff dff423(x[23],clk,reset,df4[23]);
d_ff dff424(x[24],clk,reset,df4[24]);
d_ff dff425(x[25],clk,reset,df4[25]);
d_ff dff426(x[26],clk,reset,df4[26]);
d_ff dff427(x[27],clk,reset,df4[27]);
d_ff dff428(x[28],clk,reset,df4[28]);
d_ff dff429(x[29],clk,reset,df4[29]);
d_ff dff430(x[30],clk,reset,df4[30]);
d_ff dff431(x[31],clk,reset,df4[31]);
d_ff dff432(df3[48],clk,reset,df4[32]);
d_ff dff433(df3[49],clk,reset,df4[33]);
//stage 6
dot d32(cout1,df4[32],df4[33],df4[31]);
d_ff dff500(df4[0],clk,reset,df5[0]);
d_ff dff501(df4[1],clk,reset,df5[1]);
d_ff dff502(df4[2],clk,reset,df5[2]);
d_ff dff503(df4[3],clk,reset,df5[3]);
d_ff dff504(df4[4],clk,reset,df5[4]);
d_ff dff505(df4[5],clk,reset,df5[5]);
d_ff dff506(df4[6],clk,reset,df5[6]);
d_ff dff507(df4[7],clk,reset,df5[7]);
d_ff dff508(df4[8],clk,reset,df5[8]);
d_ff dff509(df4[9],clk,reset,df5[9]);
d_ff dff510(df4[10],clk,reset,df5[10]);
d_ff dff511(df4[11],clk,reset,df5[11]);
d_ff dff512(df4[12],clk,reset,df5[12]);
d_ff dff513(df4[13],clk,reset,df5[13]);
d_ff dff514(df4[14],clk,reset,df5[14]);
d_ff dff515(df4[15],clk,reset,df5[15]);
d_ff dff516(df4[16],clk,reset,df5[16]);
d_ff dff517(df4[17],clk,reset,df5[17]);
d_ff dff518(df4[18],clk,reset,df5[18]);
d_ff dff519(df4[19],clk,reset,df5[19]);
d_ff dff520(df4[20],clk,reset,df5[20]);
d_ff dff521(df4[21],clk,reset,df5[21]);
d_ff dff522(df4[22],clk,reset,df5[22]);
d_ff dff523(df4[23],clk,reset,df5[23]);
d_ff dff524(df4[24],clk,reset,df5[24]);
d_ff dff525(df4[25],clk,reset,df5[25]);
d_ff dff526(df4[26],clk,reset,df5[26]);
d_ff dff527(df4[27],clk,reset,df5[27]);
d_ff dff528(df4[28],clk,reset,df5[28]);
d_ff dff529(df4[29],clk,reset,df5[29]);
d_ff dff530(df4[30],clk,reset,df5[30]);
d_ff dff531(df4[31],clk,reset,df5[31]);
d_ff dff532(df4[32],clk,reset,df5[32]);
d_ff dff533(df4[33],clk,reset,df5[33]);
d_ff dff534(cout1,clk,reset,cout2);
assign s=df5[31:0]^p;
assign cout=cout2;
endmodule
