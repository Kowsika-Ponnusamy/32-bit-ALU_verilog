module wallacepipe32(out,x,y,clk,reset);
input [31:0]x,y;
input clk,reset;
output [63:0] out;
wire cout,over;
wire [31:0]z0,z1,z2,z3,z4,z5,z6,z7,z8,z9,z10,z11,z12,z13,z14,z15,z16,z17,z18,z19,z20,z21,z22,z23,z24,z25,z26,z27,z28,z29,z30,z31;
wire [63:0] a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15,a16,a17,a18,a19,a20,a21,a22,a23,a24,a25,a26,a27,a28,a29,a30,a31;
wire [63:0] q0,q1,q2,q3,q4,q5,q6,q7,q8,q9,q10,q11,q12,q13,q14,q15,q16,q17,q18,q19,q20,q21,q22,q23,q24,q25,q26,q27,q28,q29,q30,q31;
wire [63:0] s0,s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,s16,s17,s18,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29;
wire [63:0] sx0,sx1,sx2,sx3,sx4,sx5,sx6,sx7,sx8,sx9,sx10,sx11,sx12,sx13,sx14,sx15,sx16,sx17,sx18,sx19,sx20,sx21,sx22,sx23,sx24,sx25,sx26,sx27,sx28,sx29;
wire [63:0] c0,c1,c2,c3,c4,c5,c6,c7,c8,c9,c10,c11,c12,c13,c14,c15,c16,c17,c18,c19,c20,c21,c22,c23,c24,c25,c26,c27,c28,c29;
wire [63:0] cx0,cx1,cx2,cx3,cx4,cx5,cx6,cx7,cx8,cx9,cx10,cx11,cx12,cx13,cx14,cx15,cx16,cx17,cx18,cx19,cx20,cx21,cx22,cx23,cx24,cx25,cx26,cx27,cx28,cx29;
wire [63:0] q130,q131,q231,q331,q431,q531,q532,q631;

assign z0[0]=x[0]&y[0];
assign z0[1]=x[1]&y[0];
assign z0[2]=x[2]&y[0];
assign z0[3]=x[3]&y[0];
assign z0[4]=x[4]&y[0];
assign z0[5]=x[5]&y[0];
assign z0[6]=x[6]&y[0];
assign z0[7]=x[7]&y[0];
assign z0[8]=x[8]&y[0];
assign z0[9]=x[9]&y[0];
assign z0[10]=x[10]&y[0];
assign z0[11]=x[11]&y[0];
assign z0[12]=x[12]&y[0];
assign z0[13]=x[13]&y[0];
assign z0[14]=x[14]&y[0];
assign z0[15]=x[15]&y[0];
assign z0[16]=x[16]&y[0];
assign z0[17]=x[17]&y[0];
assign z0[18]=x[18]&y[0];
assign z0[19]=x[19]&y[0];
assign z0[20]=x[20]&y[0];
assign z0[21]=x[21]&y[0];
assign z0[22]=x[22]&y[0];
assign z0[23]=x[23]&y[0];
assign z0[24]=x[24]&y[0];
assign z0[25]=x[25]&y[0];
assign z0[26]=x[26]&y[0];
assign z0[27]=x[27]&y[0];
assign z0[28]=x[28]&y[0];
assign z0[29]=x[29]&y[0];
assign z0[30]=x[30]&y[0];
assign z0[31]=x[31]&y[0];
	assign	a0[31:0]=z0;
	assign	a0[63:32]= 0;
assign z1[0]=x[0]&y[1];
assign z1[1]=x[1]&y[1];
assign z1[2]=x[2]&y[1];
assign z1[3]=x[3]&y[1];
assign z1[4]=x[4]&y[1];
assign z1[5]=x[5]&y[1];
assign z1[6]=x[6]&y[1];
assign z1[7]=x[7]&y[1];
assign z1[8]=x[8]&y[1];
assign z1[9]=x[9]&y[1];
assign z1[10]=x[10]&y[1];
assign z1[11]=x[11]&y[1];
assign z1[12]=x[12]&y[1];
assign z1[13]=x[13]&y[1];
assign z1[14]=x[14]&y[1];
assign z1[15]=x[15]&y[1];
assign z1[16]=x[16]&y[1];
assign z1[17]=x[17]&y[1];
assign z1[18]=x[18]&y[1];
assign z1[19]=x[19]&y[1];
assign z1[20]=x[20]&y[1];
assign z1[21]=x[21]&y[1];
assign z1[22]=x[22]&y[1];
assign z1[23]=x[23]&y[1];
assign z1[24]=x[24]&y[1];
assign z1[25]=x[25]&y[1];
assign z1[26]=x[26]&y[1];
assign z1[27]=x[27]&y[1];
assign z1[28]=x[28]&y[1];
assign z1[29]=x[29]&y[1];
assign z1[30]=x[30]&y[1];
assign z1[31]=x[31]&y[1];	
	assign	a1[0]=0;
	assign	a1[32:1] = z1;
	assign	a1[63:33]=0;
assign z2[0]=x[0]&y[2];
assign z2[1]=x[1]&y[2];
assign z2[2]=x[2]&y[2];
assign z2[3]=x[3]&y[2];
assign z2[4]=x[4]&y[2];
assign z2[5]=x[5]&y[2];
assign z2[6]=x[6]&y[2];
assign z2[7]=x[7]&y[2];
assign z2[8]=x[8]&y[2];
assign z2[9]=x[9]&y[2];
assign z2[10]=x[10]&y[2];
assign z2[11]=x[11]&y[2];
assign z2[12]=x[12]&y[2];
assign z2[13]=x[13]&y[2];
assign z2[14]=x[14]&y[2];
assign z2[15]=x[15]&y[2];
assign z2[16]=x[16]&y[2];
assign z2[17]=x[17]&y[2];
assign z2[18]=x[18]&y[2];
assign z2[19]=x[19]&y[2];
assign z2[20]=x[20]&y[2];
assign z2[21]=x[21]&y[2];
assign z2[22]=x[22]&y[2];
assign z2[23]=x[23]&y[2];
assign z2[24]=x[24]&y[2];
assign z2[25]=x[25]&y[2];
assign z2[26]=x[26]&y[2];
assign z2[27]=x[27]&y[2];
assign z2[28]=x[28]&y[2];
assign z2[29]=x[29]&y[2];
assign z2[30]=x[30]&y[2];
assign z2[31]=x[31]&y[2];
		assign a2[1:0]=0;
		assign a2[33:2]=z2;
		assign a2[63:34]=0;
assign z3[0]=x[0]&y[3];
assign z3[1]=x[1]&y[3];
assign z3[2]=x[2]&y[3];
assign z3[3]=x[3]&y[3];
assign z3[4]=x[4]&y[3];
assign z3[5]=x[5]&y[3];
assign z3[6]=x[6]&y[3];
assign z3[7]=x[7]&y[3];
assign z3[8]=x[8]&y[3];
assign z3[9]=x[9]&y[3];
assign z3[10]=x[10]&y[3];
assign z3[11]=x[11]&y[3];
assign z3[12]=x[12]&y[3];
assign z3[13]=x[13]&y[3];
assign z3[14]=x[14]&y[3];
assign z3[15]=x[15]&y[3];
assign z3[16]=x[16]&y[3];
assign z3[17]=x[17]&y[3];
assign z3[18]=x[18]&y[3];
assign z3[19]=x[19]&y[3];
assign z3[20]=x[20]&y[3];
assign z3[21]=x[21]&y[3];
assign z3[22]=x[22]&y[3];
assign z3[23]=x[23]&y[3];
assign z3[24]=x[24]&y[3];
assign z3[25]=x[25]&y[3];
assign z3[26]=x[26]&y[3];
assign z3[27]=x[27]&y[3];
assign z3[28]=x[28]&y[3];
assign z3[29]=x[29]&y[3];
assign z3[30]=x[30]&y[3];
assign z3[31]=x[31]&y[3];
		assign a3[2:0]=0;
		assign a3[34:3]=z3;
		assign a3[63:35]=0;
assign z4[0]=x[0]&y[4];
assign z4[1]=x[1]&y[4];
assign z4[2]=x[2]&y[4];
assign z4[3]=x[3]&y[4];
assign z4[4]=x[4]&y[4];
assign z4[5]=x[5]&y[4];
assign z4[6]=x[6]&y[4];
assign z4[7]=x[7]&y[4];
assign z4[8]=x[8]&y[4];
assign z4[9]=x[9]&y[4];
assign z4[10]=x[10]&y[4];
assign z4[11]=x[11]&y[4];
assign z4[12]=x[12]&y[4];
assign z4[13]=x[13]&y[4];
assign z4[14]=x[14]&y[4];
assign z4[15]=x[15]&y[4];
assign z4[16]=x[16]&y[4];
assign z4[17]=x[17]&y[4];
assign z4[18]=x[18]&y[4];
assign z4[19]=x[19]&y[4];
assign z4[20]=x[20]&y[4];
assign z4[21]=x[21]&y[4];
assign z4[22]=x[22]&y[4];
assign z4[23]=x[23]&y[4];
assign z4[24]=x[24]&y[4];
assign z4[25]=x[25]&y[4];
assign z4[26]=x[26]&y[4];
assign z4[27]=x[27]&y[4];
assign z4[28]=x[28]&y[4];
assign z4[29]=x[29]&y[4];
assign z4[30]=x[30]&y[4];
assign z4[31]=x[31]&y[4];
		assign a4[3:0]=0;
		assign a4[35:4]=z4;
		assign a4[63:36]=0;
assign z5[0]=x[0]&y[5];
assign z5[1]=x[1]&y[5];
assign z5[2]=x[2]&y[5];
assign z5[3]=x[3]&y[5];
assign z5[4]=x[4]&y[5];
assign z5[5]=x[5]&y[5];
assign z5[6]=x[6]&y[5];
assign z5[7]=x[7]&y[5];
assign z5[8]=x[8]&y[5];
assign z5[9]=x[9]&y[5];
assign z5[10]=x[10]&y[5];
assign z5[11]=x[11]&y[5];
assign z5[12]=x[12]&y[5];
assign z5[13]=x[13]&y[5];
assign z5[14]=x[14]&y[5];
assign z5[15]=x[15]&y[5];
assign z5[16]=x[16]&y[5];
assign z5[17]=x[17]&y[5];
assign z5[18]=x[18]&y[5];
assign z5[19]=x[19]&y[5];
assign z5[20]=x[20]&y[5];
assign z5[21]=x[21]&y[5];
assign z5[22]=x[22]&y[5];
assign z5[23]=x[23]&y[5];
assign z5[24]=x[24]&y[5];
assign z5[25]=x[25]&y[5];
assign z5[26]=x[26]&y[5];
assign z5[27]=x[27]&y[5];
assign z5[28]=x[28]&y[5];
assign z5[29]=x[29]&y[5];
assign z5[30]=x[30]&y[5];
assign z5[31]=x[31]&y[5];
		assign a5[4:0]=0;
		assign a5[36:5]=z5;
		assign a5[63:37]=0;
assign z6[0]=x[0]&y[6];
assign z6[1]=x[1]&y[6];
assign z6[2]=x[2]&y[6];
assign z6[3]=x[3]&y[6];
assign z6[4]=x[4]&y[6];
assign z6[5]=x[5]&y[6];
assign z6[6]=x[6]&y[6];
assign z6[7]=x[7]&y[6];
assign z6[8]=x[8]&y[6];
assign z6[9]=x[9]&y[6];
assign z6[10]=x[10]&y[6];
assign z6[11]=x[11]&y[6];
assign z6[12]=x[12]&y[6];
assign z6[13]=x[13]&y[6];
assign z6[14]=x[14]&y[6];
assign z6[15]=x[15]&y[6];
assign z6[16]=x[16]&y[6];
assign z6[17]=x[17]&y[6];
assign z6[18]=x[18]&y[6];
assign z6[19]=x[19]&y[6];
assign z6[20]=x[20]&y[6];
assign z6[21]=x[21]&y[6];
assign z6[22]=x[22]&y[6];
assign z6[23]=x[23]&y[6];
assign z6[24]=x[24]&y[6];
assign z6[25]=x[25]&y[6];
assign z6[26]=x[26]&y[6];
assign z6[27]=x[27]&y[6];
assign z6[28]=x[28]&y[6];
assign z6[29]=x[29]&y[6];
assign z6[30]=x[30]&y[6];
assign z6[31]=x[31]&y[6];
		assign a6[5:0]=0;
		assign a6[37:6]=z6;
		assign a6[63:38]=0;
assign z7[0]=x[0]&y[7];
assign z7[1]=x[1]&y[7];
assign z7[2]=x[2]&y[7];
assign z7[3]=x[3]&y[7];
assign z7[4]=x[4]&y[7];
assign z7[5]=x[5]&y[7];
assign z7[6]=x[6]&y[7];
assign z7[7]=x[7]&y[7];
assign z7[8]=x[8]&y[7];
assign z7[9]=x[9]&y[7];
assign z7[10]=x[10]&y[7];
assign z7[11]=x[11]&y[7];
assign z7[12]=x[12]&y[7];
assign z7[13]=x[13]&y[7];
assign z7[14]=x[14]&y[7];
assign z7[15]=x[15]&y[7];
assign z7[16]=x[16]&y[7];
assign z7[17]=x[17]&y[7];
assign z7[18]=x[18]&y[7];
assign z7[19]=x[19]&y[7];
assign z7[20]=x[20]&y[7];
assign z7[21]=x[21]&y[7];
assign z7[22]=x[22]&y[7];
assign z7[23]=x[23]&y[7];
assign z7[24]=x[24]&y[7];
assign z7[25]=x[25]&y[7];
assign z7[26]=x[26]&y[7];
assign z7[27]=x[27]&y[7];
assign z7[28]=x[28]&y[7];
assign z7[29]=x[29]&y[7];
assign z7[30]=x[30]&y[7];
assign z7[31]=x[31]&y[7];
		assign a7[6:0]=0;
		assign a7[38:7]=z7;
		assign a7[63:39]=0;
assign z8[0]=x[0]&y[8];
assign z8[1]=x[1]&y[8];
assign z8[2]=x[2]&y[8];
assign z8[3]=x[3]&y[8];
assign z8[4]=x[4]&y[8];
assign z8[5]=x[5]&y[8];
assign z8[6]=x[6]&y[8];
assign z8[7]=x[7]&y[8];
assign z8[8]=x[8]&y[8];
assign z8[9]=x[9]&y[8];
assign z8[10]=x[10]&y[8];
assign z8[11]=x[11]&y[8];
assign z8[12]=x[12]&y[8];
assign z8[13]=x[13]&y[8];
assign z8[14]=x[14]&y[8];
assign z8[15]=x[15]&y[8];
assign z8[16]=x[16]&y[8];
assign z8[17]=x[17]&y[8];
assign z8[18]=x[18]&y[8];
assign z8[19]=x[19]&y[8];
assign z8[20]=x[20]&y[8];
assign z8[21]=x[21]&y[8];
assign z8[22]=x[22]&y[8];
assign z8[23]=x[23]&y[8];
assign z8[24]=x[24]&y[8];
assign z8[25]=x[25]&y[8];
assign z8[26]=x[26]&y[8];
assign z8[27]=x[27]&y[8];
assign z8[28]=x[28]&y[8];
assign z8[29]=x[29]&y[8];
assign z8[30]=x[30]&y[8];
assign z8[31]=x[31]&y[8];
		assign a8[7:0]=0;
		assign a8[39:8]=z8;
		assign a8[63:40]=0;
assign z9[0]=x[0]&y[9];
assign z9[1]=x[1]&y[9];
assign z9[2]=x[2]&y[9];
assign z9[3]=x[3]&y[9];
assign z9[4]=x[4]&y[9];
assign z9[5]=x[5]&y[9];
assign z9[6]=x[6]&y[9];
assign z9[7]=x[7]&y[9];
assign z9[8]=x[8]&y[9];
assign z9[9]=x[9]&y[9];
assign z9[10]=x[10]&y[9];
assign z9[11]=x[11]&y[9];
assign z9[12]=x[12]&y[9];
assign z9[13]=x[13]&y[9];
assign z9[14]=x[14]&y[9];
assign z9[15]=x[15]&y[9];
assign z9[16]=x[16]&y[9];
assign z9[17]=x[17]&y[9];
assign z9[18]=x[18]&y[9];
assign z9[19]=x[19]&y[9];
assign z9[20]=x[20]&y[9];
assign z9[21]=x[21]&y[9];
assign z9[22]=x[22]&y[9];
assign z9[23]=x[23]&y[9];
assign z9[24]=x[24]&y[9];
assign z9[25]=x[25]&y[9];
assign z9[26]=x[26]&y[9];
assign z9[27]=x[27]&y[9];
assign z9[28]=x[28]&y[9];
assign z9[29]=x[29]&y[9];
assign z9[30]=x[30]&y[9];
assign z9[31]=x[31]&y[9];
		assign a9[8:0]=0;
		assign a9[40:9]=z9;
		assign a9[63:41]=0;
assign z10[0]=x[0]&y[10];
assign z10[1]=x[1]&y[10];
assign z10[2]=x[2]&y[10];
assign z10[3]=x[3]&y[10];
assign z10[4]=x[4]&y[10];
assign z10[5]=x[5]&y[10];
assign z10[6]=x[6]&y[10];
assign z10[7]=x[7]&y[10];
assign z10[8]=x[8]&y[10];
assign z10[9]=x[9]&y[10];
assign z10[10]=x[10]&y[10];
assign z10[11]=x[11]&y[10];
assign z10[12]=x[12]&y[10];
assign z10[13]=x[13]&y[10];
assign z10[14]=x[14]&y[10];
assign z10[15]=x[15]&y[10];
assign z10[16]=x[16]&y[10];
assign z10[17]=x[17]&y[10];
assign z10[18]=x[18]&y[10];
assign z10[19]=x[19]&y[10];
assign z10[20]=x[20]&y[10];
assign z10[21]=x[21]&y[10];
assign z10[22]=x[22]&y[10];
assign z10[23]=x[23]&y[10];
assign z10[24]=x[24]&y[10];
assign z10[25]=x[25]&y[10];
assign z10[26]=x[26]&y[10];
assign z10[27]=x[27]&y[10];
assign z10[28]=x[28]&y[10];
assign z10[29]=x[29]&y[10];
assign z10[30]=x[30]&y[10];
assign z10[31]=x[31]&y[10];
		assign a10[9:0]=0;
		assign a10[41:10]=z10;
		assign a10[63:41]=0;
assign z11[0]=x[0]&y[11];
assign z11[1]=x[1]&y[11];
assign z11[2]=x[2]&y[11];
assign z11[3]=x[3]&y[11];
assign z11[4]=x[4]&y[11];
assign z11[5]=x[5]&y[11];
assign z11[6]=x[6]&y[11];
assign z11[7]=x[7]&y[11];
assign z11[8]=x[8]&y[11];
assign z11[9]=x[9]&y[11];
assign z11[10]=x[10]&y[11];
assign z11[11]=x[11]&y[11];
assign z11[12]=x[12]&y[11];
assign z11[13]=x[13]&y[11];
assign z11[14]=x[14]&y[11];
assign z11[15]=x[15]&y[11];
assign z11[16]=x[16]&y[11];
assign z11[17]=x[17]&y[11];
assign z11[18]=x[18]&y[11];
assign z11[19]=x[19]&y[11];
assign z11[20]=x[20]&y[11];
assign z11[21]=x[21]&y[11];
assign z11[22]=x[22]&y[11];
assign z11[23]=x[23]&y[11];
assign z11[24]=x[24]&y[11];
assign z11[25]=x[25]&y[11];
assign z11[26]=x[26]&y[11];
assign z11[27]=x[27]&y[11];
assign z11[28]=x[28]&y[11];
assign z11[29]=x[29]&y[11];
assign z11[30]=x[30]&y[11];
assign z11[31]=x[31]&y[11];
		assign a11[10:0]=0;
		assign a11[42:11]=z11;
		assign a11[63:43]=0;
assign z12[0]=x[0]&y[12];
assign z12[1]=x[1]&y[12];
assign z12[2]=x[2]&y[12];
assign z12[3]=x[3]&y[12];
assign z12[4]=x[4]&y[12];
assign z12[5]=x[5]&y[12];
assign z12[6]=x[6]&y[12];
assign z12[7]=x[7]&y[12];
assign z12[8]=x[8]&y[12];
assign z12[9]=x[9]&y[12];
assign z12[10]=x[10]&y[12];
assign z12[11]=x[11]&y[12];
assign z12[12]=x[12]&y[12];
assign z12[13]=x[13]&y[12];
assign z12[14]=x[14]&y[12];
assign z12[15]=x[15]&y[12];
assign z12[16]=x[16]&y[12];
assign z12[17]=x[17]&y[12];
assign z12[18]=x[18]&y[12];
assign z12[19]=x[19]&y[12];
assign z12[20]=x[20]&y[12];
assign z12[21]=x[21]&y[12];
assign z12[22]=x[22]&y[12];
assign z12[23]=x[23]&y[12];
assign z12[24]=x[24]&y[12];
assign z12[25]=x[25]&y[12];
assign z12[26]=x[26]&y[12];
assign z12[27]=x[27]&y[12];
assign z12[28]=x[28]&y[12];
assign z12[29]=x[29]&y[12];
assign z12[30]=x[30]&y[12];
assign z12[31]=x[31]&y[12];
		assign a12[11:0]=0;
		assign a12[43:12]=z12;
		assign a12[63:44]=0;
assign z13[0]=x[0]&y[13];
assign z13[1]=x[1]&y[13];
assign z13[2]=x[2]&y[13];
assign z13[3]=x[3]&y[13];
assign z13[4]=x[4]&y[13];
assign z13[5]=x[5]&y[13];
assign z13[6]=x[6]&y[13];
assign z13[7]=x[7]&y[13];
assign z13[8]=x[8]&y[13];
assign z13[9]=x[9]&y[13];
assign z13[10]=x[10]&y[13];
assign z13[11]=x[11]&y[13];
assign z13[12]=x[12]&y[13];
assign z13[13]=x[13]&y[13];
assign z13[14]=x[14]&y[13];
assign z13[15]=x[15]&y[13];
assign z13[16]=x[16]&y[13];
assign z13[17]=x[17]&y[13];
assign z13[18]=x[18]&y[13];
assign z13[19]=x[19]&y[13];
assign z13[20]=x[20]&y[13];
assign z13[21]=x[21]&y[13];
assign z13[22]=x[22]&y[13];
assign z13[23]=x[23]&y[13];
assign z13[24]=x[24]&y[13];
assign z13[25]=x[25]&y[13];
assign z13[26]=x[26]&y[13];
assign z13[27]=x[27]&y[13];
assign z13[28]=x[28]&y[13];
assign z13[29]=x[29]&y[13];
assign z13[30]=x[30]&y[13];
assign z13[31]=x[31]&y[13];
		assign a13[12:0]=0;
		assign a13[44:13]=z13;
		assign a13[63:45]=0;
assign z14[0]=x[0]&y[14];
assign z14[1]=x[1]&y[14];
assign z14[2]=x[2]&y[14];
assign z14[3]=x[3]&y[14];
assign z14[4]=x[4]&y[14];
assign z14[5]=x[5]&y[14];
assign z14[6]=x[6]&y[14];
assign z14[7]=x[7]&y[14];
assign z14[8]=x[8]&y[14];
assign z14[9]=x[9]&y[14];
assign z14[10]=x[10]&y[14];
assign z14[11]=x[11]&y[14];
assign z14[12]=x[12]&y[14];
assign z14[13]=x[13]&y[14];
assign z14[14]=x[14]&y[14];
assign z14[15]=x[15]&y[14];
assign z14[16]=x[16]&y[14];
assign z14[17]=x[17]&y[14];
assign z14[18]=x[18]&y[14];
assign z14[19]=x[19]&y[14];
assign z14[20]=x[20]&y[14];
assign z14[21]=x[21]&y[14];
assign z14[22]=x[22]&y[14];
assign z14[23]=x[23]&y[14];
assign z14[24]=x[24]&y[14];
assign z14[25]=x[25]&y[14];
assign z14[26]=x[26]&y[14];
assign z14[27]=x[27]&y[14];
assign z14[28]=x[28]&y[14];
assign z14[29]=x[29]&y[14];
assign z14[30]=x[30]&y[14];
assign z14[31]=x[31]&y[14];
		assign a14[13:0]=0;
		assign a14[45:14]=z14;
		assign a14[63:46]=0;
assign z15[0]=x[0]&y[15];
assign z15[1]=x[1]&y[15];
assign z15[2]=x[2]&y[15];
assign z15[3]=x[3]&y[15];
assign z15[4]=x[4]&y[15];
assign z15[5]=x[5]&y[15];
assign z15[6]=x[6]&y[15];
assign z15[7]=x[7]&y[15];
assign z15[8]=x[8]&y[15];
assign z15[9]=x[9]&y[15];
assign z15[10]=x[10]&y[15];
assign z15[11]=x[11]&y[15];
assign z15[12]=x[12]&y[15];
assign z15[13]=x[13]&y[15];
assign z15[14]=x[14]&y[15];
assign z15[15]=x[15]&y[15];
assign z15[16]=x[16]&y[15];
assign z15[17]=x[17]&y[15];
assign z15[18]=x[18]&y[15];
assign z15[19]=x[19]&y[15];
assign z15[20]=x[20]&y[15];
assign z15[21]=x[21]&y[15];
assign z15[22]=x[22]&y[15];
assign z15[23]=x[23]&y[15];
assign z15[24]=x[24]&y[15];
assign z15[25]=x[25]&y[15];
assign z15[26]=x[26]&y[15];
assign z15[27]=x[27]&y[15];
assign z15[28]=x[28]&y[15];
assign z15[29]=x[29]&y[15];
assign z15[30]=x[30]&y[15];
assign z15[31]=x[31]&y[15];
		assign a15[14:0]=0;
		assign a15[46:15]=z15;
		assign a15[63:47]=0;
assign z16[0]=x[0]&y[16];
assign z16[1]=x[1]&y[16];
assign z16[2]=x[2]&y[16];
assign z16[3]=x[3]&y[16];
assign z16[4]=x[4]&y[16];
assign z16[5]=x[5]&y[16];
assign z16[6]=x[6]&y[16];
assign z16[7]=x[7]&y[16];
assign z16[8]=x[8]&y[16];
assign z16[9]=x[9]&y[16];
assign z16[10]=x[10]&y[16];
assign z16[11]=x[11]&y[16];
assign z16[12]=x[12]&y[16];
assign z16[13]=x[13]&y[16];
assign z16[14]=x[14]&y[16];
assign z16[15]=x[15]&y[16];
assign z16[16]=x[16]&y[16];
assign z16[17]=x[17]&y[16];
assign z16[18]=x[18]&y[16];
assign z16[19]=x[19]&y[16];
assign z16[20]=x[20]&y[16];
assign z16[21]=x[21]&y[16];
assign z16[22]=x[22]&y[16];
assign z16[23]=x[23]&y[16];
assign z16[24]=x[24]&y[16];
assign z16[25]=x[25]&y[16];
assign z16[26]=x[26]&y[16];
assign z16[27]=x[27]&y[16];
assign z16[28]=x[28]&y[16];
assign z16[29]=x[29]&y[16];
assign z16[30]=x[30]&y[16];
assign z16[31]=x[31]&y[16];
		assign a16[15:0]=0;
		assign a16[47:16]=z16;
		assign a16[63:48]=0;
assign z17[0]=x[0]&y[17];
assign z17[1]=x[1]&y[17];
assign z17[2]=x[2]&y[17];
assign z17[3]=x[3]&y[17];
assign z17[4]=x[4]&y[17];
assign z17[5]=x[5]&y[17];
assign z17[6]=x[6]&y[17];
assign z17[7]=x[7]&y[17];
assign z17[8]=x[8]&y[17];
assign z17[9]=x[9]&y[17];
assign z17[10]=x[10]&y[17];
assign z17[11]=x[11]&y[17];
assign z17[12]=x[12]&y[17];
assign z17[13]=x[13]&y[17];
assign z17[14]=x[14]&y[17];
assign z17[15]=x[15]&y[17];
assign z17[16]=x[16]&y[17];
assign z17[17]=x[17]&y[17];
assign z17[18]=x[18]&y[17];
assign z17[19]=x[19]&y[17];
assign z17[20]=x[20]&y[17];
assign z17[21]=x[21]&y[17];
assign z17[22]=x[22]&y[17];
assign z17[23]=x[23]&y[17];
assign z17[24]=x[24]&y[17];
assign z17[25]=x[25]&y[17];
assign z17[26]=x[26]&y[17];
assign z17[27]=x[27]&y[17];
assign z17[28]=x[28]&y[17];
assign z17[29]=x[29]&y[17];
assign z17[30]=x[30]&y[17];
assign z17[31]=x[31]&y[17];
		assign a17[16:0]=0;
		assign a17[48:17]=z17;
		assign a17[63:49]=0;
assign z18[0]=x[0]&y[18];
assign z18[1]=x[1]&y[18];
assign z18[2]=x[2]&y[18];
assign z18[3]=x[3]&y[18];
assign z18[4]=x[4]&y[18];
assign z18[5]=x[5]&y[18];
assign z18[6]=x[6]&y[18];
assign z18[7]=x[7]&y[18];
assign z18[8]=x[8]&y[18];
assign z18[9]=x[9]&y[18];
assign z18[10]=x[10]&y[18];
assign z18[11]=x[11]&y[18];
assign z18[12]=x[12]&y[18];
assign z18[13]=x[13]&y[18];
assign z18[14]=x[14]&y[18];
assign z18[15]=x[15]&y[18];
assign z18[16]=x[16]&y[18];
assign z18[17]=x[17]&y[18];
assign z18[18]=x[18]&y[18];
assign z18[19]=x[19]&y[18];
assign z18[20]=x[20]&y[18];
assign z18[21]=x[21]&y[18];
assign z18[22]=x[22]&y[18];
assign z18[23]=x[23]&y[18];
assign z18[24]=x[24]&y[18];
assign z18[25]=x[25]&y[18];
assign z18[26]=x[26]&y[18];
assign z18[27]=x[27]&y[18];
assign z18[28]=x[28]&y[18];
assign z18[29]=x[29]&y[18];
assign z18[30]=x[30]&y[18];
assign z18[31]=x[31]&y[18];
		assign a18[17:0]=0;
		assign a18[49:18]=z18;
		assign a18[63:50]=0;
assign z19[0]=x[0]&y[19];
assign z19[1]=x[1]&y[19];
assign z19[2]=x[2]&y[19];
assign z19[3]=x[3]&y[19];
assign z19[4]=x[4]&y[19];
assign z19[5]=x[5]&y[19];
assign z19[6]=x[6]&y[19];
assign z19[7]=x[7]&y[19];
assign z19[8]=x[8]&y[19];
assign z19[9]=x[9]&y[19];
assign z19[10]=x[10]&y[19];
assign z19[11]=x[11]&y[19];
assign z19[12]=x[12]&y[19];
assign z19[13]=x[13]&y[19];
assign z19[14]=x[14]&y[19];
assign z19[15]=x[15]&y[19];
assign z19[16]=x[16]&y[19];
assign z19[17]=x[17]&y[19];
assign z19[18]=x[18]&y[19];
assign z19[19]=x[19]&y[19];
assign z19[20]=x[20]&y[19];
assign z19[21]=x[21]&y[19];
assign z19[22]=x[22]&y[19];
assign z19[23]=x[23]&y[19];
assign z19[24]=x[24]&y[19];
assign z19[25]=x[25]&y[19];
assign z19[26]=x[26]&y[19];
assign z19[27]=x[27]&y[19];
assign z19[28]=x[28]&y[19];
assign z19[29]=x[29]&y[19];
assign z19[30]=x[30]&y[19];
assign z19[31]=x[31]&y[19];
		assign a19[18:0]=0;
		assign a19[50:19]=z19;
		assign a19[63:51]=0;
assign z20[0]=x[0]&y[20];
assign z20[1]=x[1]&y[20];
assign z20[2]=x[2]&y[20];
assign z20[3]=x[3]&y[20];
assign z20[4]=x[4]&y[20];
assign z20[5]=x[5]&y[20];
assign z20[6]=x[6]&y[20];
assign z20[7]=x[7]&y[20];
assign z20[8]=x[8]&y[20];
assign z20[9]=x[9]&y[20];
assign z20[10]=x[10]&y[20];
assign z20[11]=x[11]&y[20];
assign z20[12]=x[12]&y[20];
assign z20[13]=x[13]&y[20];
assign z20[14]=x[14]&y[20];
assign z20[15]=x[15]&y[20];
assign z20[16]=x[16]&y[20];
assign z20[17]=x[17]&y[20];
assign z20[18]=x[18]&y[20];
assign z20[19]=x[19]&y[20];
assign z20[20]=x[20]&y[20];
assign z20[21]=x[21]&y[20];
assign z20[22]=x[22]&y[20];
assign z20[23]=x[23]&y[20];
assign z20[24]=x[24]&y[20];
assign z20[25]=x[25]&y[20];
assign z20[26]=x[26]&y[20];
assign z20[27]=x[27]&y[20];
assign z20[28]=x[28]&y[20];
assign z20[29]=x[29]&y[20];
assign z20[30]=x[30]&y[20];
assign z20[31]=x[31]&y[20];
		assign a20[19:0]=0;
		assign a20[51:20]=z20;
		assign a20[63:52]=0;
assign z21[0]=x[0]&y[21];
assign z21[1]=x[1]&y[21];
assign z21[2]=x[2]&y[21];
assign z21[3]=x[3]&y[21];
assign z21[4]=x[4]&y[21];
assign z21[5]=x[5]&y[21];
assign z21[6]=x[6]&y[21];
assign z21[7]=x[7]&y[21];
assign z21[8]=x[8]&y[21];
assign z21[9]=x[9]&y[21];
assign z21[10]=x[10]&y[21];
assign z21[11]=x[11]&y[21];
assign z21[12]=x[12]&y[21];
assign z21[13]=x[13]&y[21];
assign z21[14]=x[14]&y[21];
assign z21[15]=x[15]&y[21];
assign z21[16]=x[16]&y[21];
assign z21[17]=x[17]&y[21];
assign z21[18]=x[18]&y[21];
assign z21[19]=x[19]&y[21];
assign z21[20]=x[20]&y[21];
assign z21[21]=x[21]&y[21];
assign z21[22]=x[22]&y[21];
assign z21[23]=x[23]&y[21];
assign z21[24]=x[24]&y[21];
assign z21[25]=x[25]&y[21];
assign z21[26]=x[26]&y[21];
assign z21[27]=x[27]&y[21];
assign z21[28]=x[28]&y[21];
assign z21[29]=x[29]&y[21];
assign z21[30]=x[30]&y[21];
assign z21[31]=x[31]&y[21];
		assign a21[20:0]=0;
		assign a21[52:21]=z21;
		assign a21[63:53]=0;
assign z22[0]=x[0]&y[22];
assign z22[1]=x[1]&y[22];
assign z22[2]=x[2]&y[22];
assign z22[3]=x[3]&y[22];
assign z22[4]=x[4]&y[22];
assign z22[5]=x[5]&y[22];
assign z22[6]=x[6]&y[22];
assign z22[7]=x[7]&y[22];
assign z22[8]=x[8]&y[22];
assign z22[9]=x[9]&y[22];
assign z22[10]=x[10]&y[22];
assign z22[11]=x[11]&y[22];
assign z22[12]=x[12]&y[22];
assign z22[13]=x[13]&y[22];
assign z22[14]=x[14]&y[22];
assign z22[15]=x[15]&y[22];
assign z22[16]=x[16]&y[22];
assign z22[17]=x[17]&y[22];
assign z22[18]=x[18]&y[22];
assign z22[19]=x[19]&y[22];
assign z22[20]=x[20]&y[22];
assign z22[21]=x[21]&y[22];
assign z22[22]=x[22]&y[22];
assign z22[23]=x[23]&y[22];
assign z22[24]=x[24]&y[22];
assign z22[25]=x[25]&y[22];
assign z22[26]=x[26]&y[22];
assign z22[27]=x[27]&y[22];
assign z22[28]=x[28]&y[22];
assign z22[29]=x[29]&y[22];
assign z22[30]=x[30]&y[22];
assign z22[31]=x[31]&y[22];
		assign a22[21:0]=0;
		assign a22[53:22]=z22;
		assign a22[63:54]=0;
assign z23[0]=x[0]&y[23];
assign z23[1]=x[1]&y[23];
assign z23[2]=x[2]&y[23];
assign z23[3]=x[3]&y[23];
assign z23[4]=x[4]&y[23];
assign z23[5]=x[5]&y[23];
assign z23[6]=x[6]&y[23];
assign z23[7]=x[7]&y[23];
assign z23[8]=x[8]&y[23];
assign z23[9]=x[9]&y[23];
assign z23[10]=x[10]&y[23];
assign z23[11]=x[11]&y[23];
assign z23[12]=x[12]&y[23];
assign z23[13]=x[13]&y[23];
assign z23[14]=x[14]&y[23];
assign z23[15]=x[15]&y[23];
assign z23[16]=x[16]&y[23];
assign z23[17]=x[17]&y[23];
assign z23[18]=x[18]&y[23];
assign z23[19]=x[19]&y[23];
assign z23[20]=x[20]&y[23];
assign z23[21]=x[21]&y[23];
assign z23[22]=x[22]&y[23];
assign z23[23]=x[23]&y[23];
assign z23[24]=x[24]&y[23];
assign z23[25]=x[25]&y[23];
assign z23[26]=x[26]&y[23];
assign z23[27]=x[27]&y[23];
assign z23[28]=x[28]&y[23];
assign z23[29]=x[29]&y[23];
assign z23[30]=x[30]&y[23];
assign z23[31]=x[31]&y[23];
		assign a23[22:0]=0;
		assign a23[54:23]=z23;
		assign a23[63:55]=0;
assign z24[0]=x[0]&y[24];
assign z24[1]=x[1]&y[24];
assign z24[2]=x[2]&y[24];
assign z24[3]=x[3]&y[24];
assign z24[4]=x[4]&y[24];
assign z24[5]=x[5]&y[24];
assign z24[6]=x[6]&y[24];
assign z24[7]=x[7]&y[24];
assign z24[8]=x[8]&y[24];
assign z24[9]=x[9]&y[24];
assign z24[10]=x[10]&y[24];
assign z24[11]=x[11]&y[24];
assign z24[12]=x[12]&y[24];
assign z24[13]=x[13]&y[24];
assign z24[14]=x[14]&y[24];
assign z24[15]=x[15]&y[24];
assign z24[16]=x[16]&y[24];
assign z24[17]=x[17]&y[24];
assign z24[18]=x[18]&y[24];
assign z24[19]=x[19]&y[24];
assign z24[20]=x[20]&y[24];
assign z24[21]=x[21]&y[24];
assign z24[22]=x[22]&y[24];
assign z24[23]=x[23]&y[24];
assign z24[24]=x[24]&y[24];
assign z24[25]=x[25]&y[24];
assign z24[26]=x[26]&y[24];
assign z24[27]=x[27]&y[24];
assign z24[28]=x[28]&y[24];
assign z24[29]=x[29]&y[24];
assign z24[30]=x[30]&y[24];
assign z24[31]=x[31]&y[24];
		assign a24[23:0]=0;
		assign a24[55:24]=z24;
		assign a24[63:56]=0;
assign z25[0]=x[0]&y[25];
assign z25[1]=x[1]&y[25];
assign z25[2]=x[2]&y[25];
assign z25[3]=x[3]&y[25];
assign z25[4]=x[4]&y[25];
assign z25[5]=x[5]&y[25];
assign z25[6]=x[6]&y[25];
assign z25[7]=x[7]&y[25];
assign z25[8]=x[8]&y[25];
assign z25[9]=x[9]&y[25];
assign z25[10]=x[10]&y[25];
assign z25[11]=x[11]&y[25];
assign z25[12]=x[12]&y[25];
assign z25[13]=x[13]&y[25];
assign z25[14]=x[14]&y[25];
assign z25[15]=x[15]&y[25];
assign z25[16]=x[16]&y[25];
assign z25[17]=x[17]&y[25];
assign z25[18]=x[18]&y[25];
assign z25[19]=x[19]&y[25];
assign z25[20]=x[20]&y[25];
assign z25[21]=x[21]&y[25];
assign z25[22]=x[22]&y[25];
assign z25[23]=x[23]&y[25];
assign z25[24]=x[24]&y[25];
assign z25[25]=x[25]&y[25];
assign z25[26]=x[26]&y[25];
assign z25[27]=x[27]&y[25];
assign z25[28]=x[28]&y[25];
assign z25[29]=x[29]&y[25];
assign z25[30]=x[30]&y[25];
assign z25[31]=x[31]&y[25];
		assign a25[24:0]=0;
		assign a25[56:25]=z25;
		assign a25[63:57]=0;
assign z26[0]=x[0]&y[26];
assign z26[1]=x[1]&y[26];
assign z26[2]=x[2]&y[26];
assign z26[3]=x[3]&y[26];
assign z26[4]=x[4]&y[26];
assign z26[5]=x[5]&y[26];
assign z26[6]=x[6]&y[26];
assign z26[7]=x[7]&y[26];
assign z26[8]=x[8]&y[26];
assign z26[9]=x[9]&y[26];
assign z26[10]=x[10]&y[26];
assign z26[11]=x[11]&y[26];
assign z26[12]=x[12]&y[26];
assign z26[13]=x[13]&y[26];
assign z26[14]=x[14]&y[26];
assign z26[15]=x[15]&y[26];
assign z26[16]=x[16]&y[26];
assign z26[17]=x[17]&y[26];
assign z26[18]=x[18]&y[26];
assign z26[19]=x[19]&y[26];
assign z26[20]=x[20]&y[26];
assign z26[21]=x[21]&y[26];
assign z26[22]=x[22]&y[26];
assign z26[23]=x[23]&y[26];
assign z26[24]=x[24]&y[26];
assign z26[25]=x[25]&y[26];
assign z26[26]=x[26]&y[26];
assign z26[27]=x[27]&y[26];
assign z26[28]=x[28]&y[26];
assign z26[29]=x[29]&y[26];
assign z26[30]=x[30]&y[26];
assign z26[31]=x[31]&y[26];
		assign a26[25:0]=0;
		assign a26[57:26]=z26;
		assign a26[63:58]=0;
assign z27[0]=x[0]&y[27];
assign z27[1]=x[1]&y[27];
assign z27[2]=x[2]&y[27];
assign z27[3]=x[3]&y[27];
assign z27[4]=x[4]&y[27];
assign z27[5]=x[5]&y[27];
assign z27[6]=x[6]&y[27];
assign z27[7]=x[7]&y[27];
assign z27[8]=x[8]&y[27];
assign z27[9]=x[9]&y[27];
assign z27[10]=x[10]&y[27];
assign z27[11]=x[11]&y[27];
assign z27[12]=x[12]&y[27];
assign z27[13]=x[13]&y[27];
assign z27[14]=x[14]&y[27];
assign z27[15]=x[15]&y[27];
assign z27[16]=x[16]&y[27];
assign z27[17]=x[17]&y[27];
assign z27[18]=x[18]&y[27];
assign z27[19]=x[19]&y[27];
assign z27[20]=x[20]&y[27];
assign z27[21]=x[21]&y[27];
assign z27[22]=x[22]&y[27];
assign z27[23]=x[23]&y[27];
assign z27[24]=x[24]&y[27];
assign z27[25]=x[25]&y[27];
assign z27[26]=x[26]&y[27];
assign z27[27]=x[27]&y[27];
assign z27[28]=x[28]&y[27];
assign z27[29]=x[29]&y[27];
assign z27[30]=x[30]&y[27];
assign z27[31]=x[31]&y[27];
		assign a27[26:0]=0;
		assign a27[58:27]=z27;
		assign a27[63:59]=0;
assign z28[0]=x[0]&y[28];
assign z28[1]=x[1]&y[28];
assign z28[2]=x[2]&y[28];
assign z28[3]=x[3]&y[28];
assign z28[4]=x[4]&y[28];
assign z28[5]=x[5]&y[28];
assign z28[6]=x[6]&y[28];
assign z28[7]=x[7]&y[28];
assign z28[8]=x[8]&y[28];
assign z28[9]=x[9]&y[28];
assign z28[10]=x[10]&y[28];
assign z28[11]=x[11]&y[28];
assign z28[12]=x[12]&y[28];
assign z28[13]=x[13]&y[28];
assign z28[14]=x[14]&y[28];
assign z28[15]=x[15]&y[28];
assign z28[16]=x[16]&y[28];
assign z28[17]=x[17]&y[28];
assign z28[18]=x[18]&y[28];
assign z28[19]=x[19]&y[28];
assign z28[20]=x[20]&y[28];
assign z28[21]=x[21]&y[28];
assign z28[22]=x[22]&y[28];
assign z28[23]=x[23]&y[28];
assign z28[24]=x[24]&y[28];
assign z28[25]=x[25]&y[28];
assign z28[26]=x[26]&y[28];
assign z28[27]=x[27]&y[28];
assign z28[28]=x[28]&y[28];
assign z28[29]=x[29]&y[28];
assign z28[30]=x[30]&y[28];
assign z28[31]=x[31]&y[28];
		assign a28[27:0]=0;
		assign a28[59:28]=z28;
		assign a28[63:60]=0;
assign z29[0]=x[0]&y[29];
assign z29[1]=x[1]&y[29];
assign z29[2]=x[2]&y[29];
assign z29[3]=x[3]&y[29];
assign z29[4]=x[4]&y[29];
assign z29[5]=x[5]&y[29];
assign z29[6]=x[6]&y[29];
assign z29[7]=x[7]&y[29];
assign z29[8]=x[8]&y[29];
assign z29[9]=x[9]&y[29];
assign z29[10]=x[10]&y[29];
assign z29[11]=x[11]&y[29];
assign z29[12]=x[12]&y[29];
assign z29[13]=x[13]&y[29];
assign z29[14]=x[14]&y[29];
assign z29[15]=x[15]&y[29];
assign z29[16]=x[16]&y[29];
assign z29[17]=x[17]&y[29];
assign z29[18]=x[18]&y[29];
assign z29[19]=x[19]&y[29];
assign z29[20]=x[20]&y[29];
assign z29[21]=x[21]&y[29];
assign z29[22]=x[22]&y[29];
assign z29[23]=x[23]&y[29];
assign z29[24]=x[24]&y[29];
assign z29[25]=x[25]&y[29];
assign z29[26]=x[26]&y[29];
assign z29[27]=x[27]&y[29];
assign z29[28]=x[28]&y[29];
assign z29[29]=x[29]&y[29];
assign z29[30]=x[30]&y[29];
assign z29[31]=x[31]&y[29];
		assign a29[28:0]=0;
		assign a29[60:29]=z29;
		assign a29[63:61]=0;
assign z30[0]=x[0]&y[30];
assign z30[1]=x[1]&y[30];
assign z30[2]=x[2]&y[30];
assign z30[3]=x[3]&y[30];
assign z30[4]=x[4]&y[30];
assign z30[5]=x[5]&y[30];
assign z30[6]=x[6]&y[30];
assign z30[7]=x[7]&y[30];
assign z30[8]=x[8]&y[30];
assign z30[9]=x[9]&y[30];
assign z30[10]=x[10]&y[30];
assign z30[11]=x[11]&y[30];
assign z30[12]=x[12]&y[30];
assign z30[13]=x[13]&y[30];
assign z30[14]=x[14]&y[30];
assign z30[15]=x[15]&y[30];
assign z30[16]=x[16]&y[30];
assign z30[17]=x[17]&y[30];
assign z30[18]=x[18]&y[30];
assign z30[19]=x[19]&y[30];
assign z30[20]=x[20]&y[30];
assign z30[21]=x[21]&y[30];
assign z30[22]=x[22]&y[30];
assign z30[23]=x[23]&y[30];
assign z30[24]=x[24]&y[30];
assign z30[25]=x[25]&y[30];
assign z30[26]=x[26]&y[30];
assign z30[27]=x[27]&y[30];
assign z30[28]=x[28]&y[30];
assign z30[29]=x[29]&y[30];
assign z30[30]=x[30]&y[30];
assign z30[31]=x[31]&y[30];
		assign a30[29:0]=0;
		assign a30[61:30]=z30;
		assign a30[63:62]=0;
assign z31[0]=x[0]&y[31];
assign z31[1]=x[1]&y[31];
assign z31[2]=x[2]&y[31];
assign z31[3]=x[3]&y[31];
assign z31[4]=x[4]&y[31];
assign z31[5]=x[5]&y[31];
assign z31[6]=x[6]&y[31];
assign z31[7]=x[7]&y[31];
assign z31[8]=x[8]&y[31];
assign z31[9]=x[9]&y[31];
assign z31[10]=x[10]&y[31];
assign z31[11]=x[11]&y[31];
assign z31[12]=x[12]&y[31];
assign z31[13]=x[13]&y[31];
assign z31[14]=x[14]&y[31];
assign z31[15]=x[15]&y[31];
assign z31[16]=x[16]&y[31];
assign z31[17]=x[17]&y[31];
assign z31[18]=x[18]&y[31];
assign z31[19]=x[19]&y[31];
assign z31[20]=x[20]&y[31];
assign z31[21]=x[21]&y[31];
assign z31[22]=x[22]&y[31];
assign z31[23]=x[23]&y[31];
assign z31[24]=x[24]&y[31];
assign z31[25]=x[25]&y[31];
assign z31[26]=x[26]&y[31];
assign z31[27]=x[27]&y[31];
assign z31[28]=x[28]&y[31];
assign z31[29]=x[29]&y[31];
assign z31[30]=x[30]&y[31];
assign z31[31]=x[31]&y[31];
		assign a31[30:0]=0;
		assign a31[62:31]=z31;
		assign a31[63]=0;

dff63 df0(a0,clk,reset,q0);
dff63 df1(a1,clk,reset,q1);
dff63 df2(a2,clk,reset,q2);
dff63 df3(a3,clk,reset,q3);
dff63 df4(a4,clk,reset,q4);
dff63 df5(a5,clk,reset,q5);
dff63 df6(a6,clk,reset,q6);
dff63 df7(a7,clk,reset,q7);
dff63 df8(a8,clk,reset,q8);
dff63 df9(a9,clk,reset,q9);
dff63 df10(a10,clk,reset,q10);
dff63 df11(a11,clk,reset,q11);
dff63 df12(a12,clk,reset,q12);
dff63 df13(a13,clk,reset,q13);
dff63 df14(a14,clk,reset,q14);
dff63 df15(a15,clk,reset,q15);
dff63 df16(a16,clk,reset,q16);
dff63 df17(a17,clk,reset,q17);
dff63 df18(a18,clk,reset,q18);
dff63 df19(a19,clk,reset,q19);
dff63 df20(a20,clk,reset,q20);
dff63 df21(a21,clk,reset,q21);
dff63 df22(a22,clk,reset,q22);
dff63 df23(a23,clk,reset,q23);
dff63 df24(a24,clk,reset,q24);
dff63 df25(a25,clk,reset,q25);
dff63 df26(a26,clk,reset,q26);
dff63 df27(a27,clk,reset,q27);
dff63 df28(a28,clk,reset,q28);
dff63 df29(a29,clk,reset,q29);
dff63 df30(a30,clk,reset,q30);
dff63 df31(a31,clk,reset,q31);

csa cs0(s0,c0,q0,q1,q2);
csa cs1(s1,c1,q3,q4,q5);
csa cs2(s2,c2,q6,q7,q8);
csa cs3(s3,c3,q9,q10,q11);
csa cs4(s4,c4,q12,q13,q14);
csa cs5(s5,c5,q15,q16,q17);
csa cs6(s6,c6,q18,q19,q20);
csa cs7(s7,c7,q21,q22,q23);
csa cs8(s8,c8,q24,q25,q26);
csa cs9(s9,c9,q27,q28,q29);
dff63 df110(s0,clk,reset,sx0);
dff63 df111(s1,clk,reset,sx1);
dff63 df112(s2,clk,reset,sx2);
dff63 df113(s3,clk,reset,sx3);
dff63 df114(s4,clk,reset,sx4);
dff63 df115(s5,clk,reset,sx5);
dff63 df116(s6,clk,reset,sx6);
dff63 df117(s7,clk,reset,sx7);
dff63 df118(s8,clk,reset,sx8);
dff63 df119(s9,clk,reset,sx9);
dff63 df120(c0,clk,reset,cx0);
dff63 df121(c1,clk,reset,cx1);
dff63 df122(c2,clk,reset,cx2);
dff63 df123(c3,clk,reset,cx3);
dff63 df124(c4,clk,reset,cx4);
dff63 df125(c5,clk,reset,cx5);
dff63 df126(c6,clk,reset,cx6);
dff63 df127(c7,clk,reset,cx7);
dff63 df128(c8,clk,reset,cx8);
dff63 df129(c9,clk,reset,cx9);
dff63 df1130(q30,clk,reset,q130);
dff63 df1131(q31,clk,reset,q131);

csa cs10(s10,c10,sx0,cx0,sx1);
csa cs11(s11,c11,cx1,sx2,cx2);
csa cs12(s12,c12,sx3,cx3,sx4);
csa cs13(s13,c13,cx4,sx5,cx5);
csa cs14(s14,c14,sx6,cx6,sx7);
csa cs15(s15,c15,cx7,sx8,cx8);
csa cs16(s16,c16,sx9,cx9,q130);
dff63 df210(s10,clk,reset,sx10);
dff63 df211(s11,clk,reset,sx11);
dff63 df212(s12,clk,reset,sx12);
dff63 df213(s13,clk,reset,sx13);
dff63 df214(s14,clk,reset,sx14);
dff63 df215(s15,clk,reset,sx15);
dff63 df216(s16,clk,reset,sx16);
dff63 df220(c10,clk,reset,cx10);
dff63 df221(c11,clk,reset,cx11);
dff63 df222(c12,clk,reset,cx12);
dff63 df223(c13,clk,reset,cx13);
dff63 df224(c14,clk,reset,cx14);
dff63 df225(c15,clk,reset,cx15);
dff63 df226(c16,clk,reset,cx16);
dff63 df2131(q131,clk,reset,q231);

csa cs17(s17,c17,sx10,cx10,sx11);
csa cs18(s18,c18,cx11,sx12,cx12);
csa cs19(s19,c19,sx13,cx13,sx14);
csa cs20(s20,c20,cx14,sx15,cx15);
csa cs21(s21,c21,sx16,cx16,q231);
dff63 df310(s17,clk,reset,sx17);
dff63 df311(s18,clk,reset,sx18);
dff63 df312(s19,clk,reset,sx19);
dff63 df313(s20,clk,reset,sx20);
dff63 df314(s21,clk,reset,sx21);
dff63 df320(c17,clk,reset,cx17);
dff63 df321(c18,clk,reset,cx18);
dff63 df322(c19,clk,reset,cx19);
dff63 df323(c20,clk,reset,cx20);
dff63 df324(c21,clk,reset,cx21);


csa cs22(s22,c22,sx17,cx17,sx18);
csa cs23(s23,c23,cx18,sx19,cx19);
csa cs24(s24,c24,sx20,cx20,sx21);
dff63 df410(s22,clk,reset,sx22);
dff63 df411(s23,clk,reset,sx23);
dff63 df412(s24,clk,reset,sx24);
dff63 df420(c22,clk,reset,cx22);
dff63 df421(c23,clk,reset,cx23);
dff63 df422(c24,clk,reset,cx24);
dff63 df4131(cx21,clk,reset,q331);

csa cs25(s25,c25,sx22,cx22,sx23);
csa cs26(s26,c26,cx23,sx24,cx24);
dff63 df510(s25,clk,reset,sx25);
dff63 df511(s26,clk,reset,sx26);
dff63 df520(c25,clk,reset,cx25);
dff63 df521(c26,clk,reset,cx26);
dff63 df5131(q331,clk,reset,q431);

csa cs27(s27,c27,sx25,cx25,sx26);
dff63 df610(s27,clk,reset,sx27);
dff63 df620(c27,clk,reset,cx27);
dff63 df6131(q431,clk,reset,q531);
dff63 df6132(cx26,clk,reset,q532);

csa cs28(s28,c28,sx27,cx27,q532);
dff63 df710(s28,clk,reset,sx28);
dff63 df720(c28,clk,reset,cx28);
dff63 df7131(q531,clk,reset,q631);

csa cs29(s29,c29,sx28,cx28,q631);
dff63 df810(s29,clk,reset,sx29);
dff63 df820(c29,clk,reset,cx29);


prefix32pipe p1(out[31:0],over,sx29[31:0],cx29[31:0],0,clk,reset);
prefix32pipe p2(out[63:32],cout,sx29[63:32],cx29[63:32],over,clk,reset);
endmodule
