module prefix32(s,cout,a,b,c);
input [31:0] a,b;
input c;
output[31:0] s;
output cout;
wire [31:0]p,g,k;
wire [31:0]x;
assign p=a^b;
assign g=a&b;
assign k=g|p;
wire g12,g34,g56,g78,g910,g1112,g1314,g1516,g1718,g1920,g2122,g2324,g2526,g2728,g2930,g35,g36,g79,g710,g711,g712,g713,g714,g1113,g1114,g1921,g1922,g2325,g2326,g2729,g2730;
wire k12,k34,k56,k78,k910,k1112,k1314,k1516,k1718,k1920,k2122,k2324,k2526,k2728,k2930,k35,k36,k79,k710,k711,k712,k713,k714,k1113,k1114,k1921,k1922,k2325,k2326,k2729,k2730;
wire g1517,g1518,g1519,g1520,g1521,g1522,g1523,g1524,g1525,g1526,g1527,g1528,g1529,g1530,g2327,g2328,g2329,g2330;
wire k1517,k1518,k1519,k1520,k1521,k1522,k1523,k1534,k1525,k1526,k1527,k1528,k1529,k1530,k2327,k2328,k2329,k2330;
assign x[0]=c;

dot d1(x[1],g[0],k[0],x[0]);
circle c1(g[2],k[2],g[1],k[1],g12,k12);
circle c2(g[4],k[4],g[3],k[3],g34,k34);
circle c3(g[6],k[6],g[5],k[5],g56,k56);
circle c4(g[8],k[8],g[7],k[7],g78,k78);
circle c5(g[10],k[10],g[9],k[9],g910,k910);
circle c6(g[12],k[12],g[11],k[11],g1112,k1112);
circle c7(g[14],k[14],g[13],k[13],g1314,k1314);
circle c8(g[16],k[16],g[15],k[15],g1516,k1516);
circle c9(g[18],k[18],g[17],k[17],g1718,k1718);
circle c10(g[20],k[20],g[19],k[19],g1920,k1920);
circle c11(g[22],k[22],g[21],k[21],g2122,k2122);
circle c12(g[24],k[24],g[23],k[23],g2324,k2324);
circle c13(g[26],k[26],g[25],k[25],g2526,k2526);
circle c14(g[28],k[28],g[27],k[27],g2728,k2728);
circle c15(g[30],k[30],g[29],k[29],g2930,k2930);


dot d2(x[2],g[1],k[1],x[1]);
dot d3(x[3],g12,k12,x[1]);
circle c16(g[5],k[5],g34,k34,g35,k35);
circle c17(g56,k56,g34,k34,g36,k36);
circle c18(g[9],k[9],g78,k78,g79,k79);
circle c19(g910,k910,g78,k78,g710,k710);
circle c20(g[13],k[13],g1112,k1112,g1113,k1113);
circle c21(g1314,k1314,g1112,k1112,g1114,k1114);
circle c22(g[17],k[17],g1516,k1516,g1517,k1517);
circle c23(g1718,k1718,g1516,k1516,g1518,k1518);
circle c24(g[21],k[21],g1920,k1920,g1921,k1921);
circle c25(g2122,k2122,g1920,k1920,g1922,k1922);
circle c26(g[25],k[25],g2324,k2324,g2325,k2325);
circle c27(g2526,k2526,g2324,k2324,g2326,k2326);
circle c28(g[29],k[29],g2728,k2728,g2729,k2729);
circle c29(g2930,k2930,g2728,k2728,g2730,k2730);


dot d4(x[4],g[3],k[3],x[3]);
dot d5(x[5],g34,k34,x[3]);
dot d6(x[6],g35,k35,x[3]);
dot d7(x[7],g36,k36,x[3]);
circle c30(g[11],k[11],g710,k710,g711,k711);
circle c31(g1112,k1112,g710,k710,g712,k712);
circle c32(g1113,k1113,g710,k710,g713,k713);
circle c33(g1114,k1114,g710,k710,g714,k714);
circle c34(g[19],k[19],g1518,k1518,g1519,k1519);
circle c35(g1920,k1920,g1518,k1518,g1520,k1520);
circle c36(g1921,k1921,g1518,k1518,g1521,k1521);
circle c37(g1922,k1922,g1518,k1518,g1522,k1522);
circle c38(g[27],k[27],g2326,k2326,g2327,k2327);
circle c39(g2728,k2728,g2326,k2326,g2328,k2328);
circle c40(g2729,k2729,g2326,k2326,g2329,k2329);
circle c41(g2730,k2730,g2326,k2326,g2330,k2330);

dot d8(x[8],g[7],k[7],x[7]);
dot d9(x[9],g78,k78,x[7]);
dot d10(x[10],g79,k79,x[7]);
dot d11(x[11],g710,k710,x[7]);
dot d12(x[12],g711,k711,x[7]);
dot d13(x[13],g712,k712,x[7]);
dot d14(x[14],g713,k713,x[7]);
dot d15(x[15],g714,k714,x[7]);
circle c42(g[23],k[23],g1522,k1522,g1523,k1523);
circle c43(g2324,k2324,g1522,k1522,g1524,k1524);
circle c44(g2325,k2325,g1522,k1522,g1525,k1525);
circle c45(g2326,k2326,g1522,k1522,g1526,k1526);
circle c46(g2327,k2327,g1522,k1522,g1527,k1527);
circle c47(g2328,k2328,g1522,k1522,g1528,k1528);
circle c48(g2329,k2329,g1522,k1522,g1529,k1529);
circle c49(g2330,k2330,g1522,k1522,g1530,k1530);

dot d16(x[16],g[15],k[15],x[15]);
dot d17(x[17],g1516,k1516,x[15]);
dot d18(x[18],g1517,k1517,x[15]);
dot d19(x[19],g1518,k1518,x[15]);
dot d20(x[20],g1519,k1519,x[15]);
dot d21(x[21],g1520,k1520,x[15]);
dot d22(x[22],g1521,k1521,x[15]);
dot d23(x[23],g1522,k1522,x[15]);
dot d24(x[24],g1523,k1523,x[15]);
dot d25(x[25],g1524,k1524,x[15]);
dot d26(x[26],g1525,k1525,x[15]);
dot d27(x[27],g1526,k1526,x[15]);
dot d28(x[28],g1527,k1527,x[15]);
dot d29(x[29],g1528,k1528,x[15]);
dot d30(x[30],g1529,k1529,x[15]);
dot d31(x[31],g1530,k1530,x[15]);
dot d32(cout,g[31],k[31],x[31]);
assign s=x^p;
endmodule
